* C:\Users\alexm\Documents\1rUAB\EE\Practica3\ejercicio3\Schematic.sch

* Schematics Version 9.1 - Web Update 1
* Tue Oct 29 18:18:22 2024



** Analysis setup **
.tran 0m 3m
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic.net"
.INC "Schematic.als"


.probe


.END
