* C:\Users\Alex\Documents\1rUAB\EE\Practica3\ejercicio4\Schematic2.sch

* Schematics Version 9.1 - Web Update 1
* Tue Oct 29 12:20:52 2024



** Analysis setup **
.ac DEC 10 0.01 1.0K
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic2.net"
.INC "Schematic2.als"


.probe


.END
