* C:\Users\alexm\Documents\1rUAB\EE\Practica3\ejercicio5\Schematic2.sch

* Schematics Version 9.1 - Web Update 1
* Tue Oct 29 18:55:52 2024



** Analysis setup **
.tran 0m 0.4m
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic2.net"
.INC "Schematic2.als"


.probe


.END
